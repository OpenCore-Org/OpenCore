package ds_op_pkg;

    localparam DS_WRITE_B32 = 8'd13;
    localparam DS_WRITE2_B32 = 8'd14;

    localparam DS_READ_B32 = 8'd54;
    localparam DS_READ2_B32 = 8'd55;
endpackage
