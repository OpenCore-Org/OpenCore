`timescale 1ps/1ps


package common_pkg;

localparam THREADS_PER_WAVEFRONT = 32;
localparam MAX_WAVEFRONT_CNT = 4;
localparam WAVEFRONT_WIDTH = $clog2(MAX_WAVEFRONT_CNT);

// Number of intermediated registers between EX1
localparam SSRC_REG_CNT = 4;
localparam VSRC_REG_CNT = 8;

// Scalar enums/typedefs
typedef enum logic [2:0] {
    SOP2,
    SOP1,
    SOPK,
    SOPP,
    SOPC
} scalar_inst_format_e;

typedef struct packed {
    scalar_inst_format_e format;
    logic [7:0]  op;
    logic [7:0]  src0;
    logic [7:0]  src1;
    logic [6:0]  dst;
    logic [15:0] imm16;
    logic [31:0] literal;
} scalar_inst_t;

// Vector enums/typedefs
typedef enum logic [2:0] {
    VOP2,
    VOP1,
    VOPC,
    VINTRP,
    VOP3,
    VOP3P
} vector_inst_format_e;

typedef struct packed {
    logic [2:0] lane_sel0;
    logic [2:0] lane_sel1;
    logic [2:0] lane_sel2;
    logic [2:0] lane_sel3;
    logic [2:0] lane_sel4;
    logic [2:0] lane_sel5;
    logic [2:0] lane_sel6;
    logic [2:0] lane_sel7;
} vector_inst_dpp8_t;

typedef struct packed {
    logic [8:0] dpp_ctrl;
    logic       fi;
    logic       bc;
    logic       src0_neg;
    logic       src0_abs;
    logic       src1_neg;
    logic       src1_abs;
    logic [3:0] bank_mask;
    logic [3:0] row_mask;
} vector_inst_dpp16_t;

typedef struct packed {
    logic [7:0] src0;
    vector_inst_dpp16_t dpp16;
    vector_inst_dpp8_t dpp8;
} vector_inst_dpp_t;

typedef struct packed {
    logic [7:0] src0;
    logic [6:0] sdst;
    logic       sd;
    logic [2:0] dst_sel;
    logic [1:0] dst_u;
    logic       clmp;
    logic [1:0] omod;
    logic [2:0] src0_sel;
    logic       src0_sext;
    logic       src0_neg;
    logic       src0_abs;
    logic       s0;
    logic [2:0] src1_sel;
    logic       src1_sext;
    logic       src1_neg;
    logic       src1_abs;
    logic       s1;
} vector_inst_sdwa_t;

typedef struct packed {
    vector_inst_format_e format;
    logic [9:0] op;
    logic [8:0] src0;
    logic [8:0] src1; // Also used as VSRC1 for relevant instructions
    logic [8:0] src2;
    logic [7:0] vdst;
    logic [6:0] sdst; // Only used as SDST for VOP3B
    logic [5:0] attr;
    logic [1:0] attr_chan;
    logic       clmp;
    logic [3:0] op_sel;
    logic [2:0] op_sel_hi;
    logic [2:0] abs;
    logic [2:0] neg;
    logic [2:0] neg_hi;
    logic [1:0] omod;
    logic [31:0] literal;
    vector_inst_sdwa_t sdwa;
    vector_inst_dpp_t dpp;
} vector_inst_t;

// Flat typedefs
typedef struct packed {
    logic [11:0] offset;
    logic        dlc;
    logic        lds;
    logic [1:0]  seg;
    logic        glc;
    logic        slc;
    logic [6:0]  op;
    logic [7:0]  addr;
    logic [7:0]  data;
    logic [6:0]  saddr;
    logic [7:0]  vdst;
} flat_inst_t;

// Datashare typedefs
typedef struct packed {
    logic [7:0] offset0;
    logic [7:0] offset1;
    logic       gds;
    logic [7:0] op;
    logic [7:0] addr;
    logic [7:0] data0;
    logic [7:0] data1;
    logic [7:0] vdst;
} ds_inst_t;

// Export tyepdefs
typedef struct packed {
    logic [3:0] en;
    logic [5:0] target;
    logic       compr;
    logic       done;
    logic       vm;
    logic [7:0] vsrc0;
    logic [7:0] vsrc1;
    logic [7:0] vsrc2;
    logic [7:0] vsrc3;
} export_inst_t;

// Vector Memory Image Format
typedef struct packed {
    logic [1:0] nsa;
    logic [2:0] dim;
    logic       dlc;
    logic [3:0] dmask;
    logic       unrm;
    logic       glc;
    logic       r128;
    logic       tfe;
    logic       lwe;
    logic [7:0] op;
    logic       slc;
    logic [7:0] vaddr;
    logic [7:0] vdata;
    logic [4:0] srsrc;
    logic [4:0] ssamp;
    logic       a16;
    logic       d16;
    logic [7:0] addr1;
    logic [7:0] addr2;
    logic [7:0] addr3;
    logic [7:0] addr4;
    logic [7:0] addr5;
    logic [7:0] addr6;
    logic [7:0] addr7;
    logic [7:0] addr8;
    logic [7:0] addr9;
    logic [7:0] addr10;
    logic [7:0] addr11;
    logic [7:0] addr12;
} mimg_inst_t;

// Vector Memory Buffer Format 
typedef enum logic {
    MTBUF,
    MUBUF
} mbuf_inst_type_e;

typedef struct packed {
    mbuf_inst_type_e mbuf_type;
    logic [11:0] offset;
    logic        offen;
    logic        idxen;
    logic        glc;
    logic        dlc;
    logic        lds; // MUBUF Specific
    logic [7:0]  op; // MUBUF 8 bits vs MTBUF 4 bits
    logic [6:0]  dfmt; // MTBUF Specific
    logic [7:0]  vaddr;
    logic [7:0]  vdata;
    logic [4:0]  srsrc;
    logic        tfe;
    logic        slc;
    logic [7:0]  soffset;
} mbuf_inst_t;

typedef struct packed {
    logic [5:0]  sbase;
    logic [6:0]  sdata;
    logic        dlc;
    logic        glc;
    logic [7:0]  op;
    logic [20:0] offset; // Refers to SIGNED offset
    logic [6:0] soffset; // Strangely refers to SGPR which supplies an UNSIGNED byte offset 
} smem_inst_t;

// Common Defines 
`define FP32_0_5 32'h3F000000
`define FP32_NEG_0_5 32'hBF000000
`define FP32_1_0 32'h3F800000
`define FP32_NEG_1_0 32'hBF800000
`define FP32_2_0 32'h40000000
`define FP32_NEG_2_0 32'hC0000000
`define FP32_4_0 32'h40800000
`define FP32_NEG_4_0 32'hC0800000
`define FP32_INV_2_PI 32'h3E22F983


// Scalar Source Localparams
localparam SGPR0 = 8'd0;
localparam SGPR1 = 8'd1;
localparam SGPR2 = 8'd2;
localparam SGPR3 = 8'd3;
localparam SGPR4 = 8'd4;
localparam SGPR5 = 8'd5;
localparam SGPR6 = 8'd6;
localparam SGPR7 = 8'd7;
localparam SGPR8 = 8'd8;
localparam SGPR9 = 8'd9;
localparam SGPR10 = 8'd10;
localparam SGPR11 = 8'd11;
localparam SGPR12 = 8'd12;
localparam SGPR13 = 8'd13;
localparam SGPR14 = 8'd14;
localparam SGPR15 = 8'd15;
localparam SGPR16 = 8'd16;
localparam SGPR17 = 8'd17;
localparam SGPR18 = 8'd18;
localparam SGPR19 = 8'd19;
localparam SGPR20 = 8'd20;
localparam SGPR21 = 8'd21;
localparam SGPR22 = 8'd22;
localparam SGPR23 = 8'd23;
localparam SGPR24 = 8'd24;
localparam SGPR25 = 8'd25;
localparam SGPR26 = 8'd26;
localparam SGPR27 = 8'd27;
localparam SGPR28 = 8'd28;
localparam SGPR29 = 8'd29;
localparam SGPR30 = 8'd30;
localparam SGPR31 = 8'd31;
localparam SGPR32 = 8'd32;
localparam SGPR33 = 8'd33;
localparam SGPR34 = 8'd34;
localparam SGPR35 = 8'd35;
localparam SGPR36 = 8'd36;
localparam SGPR37 = 8'd37;
localparam SGPR38 = 8'd38;
localparam SGPR39 = 8'd39;
localparam SGPR40 = 8'd40;
localparam SGPR41 = 8'd41;
localparam SGPR42 = 8'd42;
localparam SGPR43 = 8'd43;
localparam SGPR44 = 8'd44;
localparam SGPR45 = 8'd45;
localparam SGPR46 = 8'd46;
localparam SGPR47 = 8'd47;
localparam SGPR48 = 8'd48;
localparam SGPR49 = 8'd49;
localparam SGPR50 = 8'd50;
localparam SGPR51 = 8'd51;
localparam SGPR52 = 8'd52;
localparam SGPR53 = 8'd53;
localparam SGPR54 = 8'd54;
localparam SGPR55 = 8'd55;
localparam SGPR56 = 8'd56;
localparam SGPR57 = 8'd57;
localparam SGPR58 = 8'd58;
localparam SGPR59 = 8'd59;
localparam SGPR60 = 8'd60;
localparam SGPR61 = 8'd61;
localparam SGPR62 = 8'd62;
localparam SGPR63 = 8'd63;
localparam SGPR64 = 8'd64;
localparam SGPR65 = 8'd65;
localparam SGPR66 = 8'd66;
localparam SGPR67 = 8'd67;
localparam SGPR68 = 8'd68;
localparam SGPR69 = 8'd69;
localparam SGPR70 = 8'd70;
localparam SGPR71 = 8'd71;
localparam SGPR72 = 8'd72;
localparam SGPR73 = 8'd73;
localparam SGPR74 = 8'd74;
localparam SGPR75 = 8'd75;
localparam SGPR76 = 8'd76;
localparam SGPR77 = 8'd77;
localparam SGPR78 = 8'd78;
localparam SGPR79 = 8'd79;
localparam SGPR80 = 8'd80;
localparam SGPR81 = 8'd81;
localparam SGPR82 = 8'd82;
localparam SGPR83 = 8'd83;
localparam SGPR84 = 8'd84;
localparam SGPR85 = 8'd85;
localparam SGPR86 = 8'd86;
localparam SGPR87 = 8'd87;
localparam SGPR88 = 8'd88;
localparam SGPR89 = 8'd89;
localparam SGPR90 = 8'd90;
localparam SGPR91 = 8'd91;
localparam SGPR92 = 8'd92;
localparam SGPR93 = 8'd93;
localparam SGPR94 = 8'd94;
localparam SGPR95 = 8'd95;
localparam SGPR96 = 8'd96;
localparam SGPR97 = 8'd97;
localparam SGPR98 = 8'd98;
localparam SGPR99 = 8'd99;
localparam SGPR100 = 8'd100;
localparam SGPR101 = 8'd101;
localparam SGPR102 = 8'd102;
localparam SGPR103 = 8'd103;
localparam SGPR104 = 8'd104;
localparam SGPR105 = 8'd105;

// Other values
localparam VCC_LO = 8'd106;
localparam VCC_HI = 8'd107;

// TTMP0 to TTMP15
localparam TTMP0 = 8'd108;
localparam TTMP1 = 8'd109;
localparam TTMP2 = 8'd110;
localparam TTMP3 = 8'd111;
localparam TTMP4 = 8'd112;
localparam TTMP5 = 8'd113;
localparam TTMP6 = 8'd114;
localparam TTMP7 = 8'd115;
localparam TTMP8 = 8'd116;
localparam TTMP9 = 8'd117;
localparam TTMP10 = 8'd118;
localparam TTMP11 = 8'd119;
localparam TTMP12 = 8'd120;
localparam TTMP13 = 8'd121;
localparam TTMP14 = 8'd122;
localparam TTMP15 = 8'd123;

// Other values
localparam M0 = 8'd124;
localparam NULL_ADDR = 8'd125;
localparam EXEC_LO = 8'd126;
localparam EXEC_HI = 8'd127;
localparam ZERO = 8'd128;

// INT1 to INT64
localparam INT1 = 8'd129;
localparam INT2 = 8'd130;
localparam INT3 = 8'd131;
localparam INT4 = 8'd132;
localparam INT5 = 8'd133;
localparam INT6 = 8'd134;
localparam INT7 = 8'd135;
localparam INT8 = 8'd136;
localparam INT9 = 8'd137;
localparam INT10 = 8'd138;
localparam INT11 = 8'd139;
localparam INT12 = 8'd140;
localparam INT13 = 8'd141;
localparam INT14 = 8'd142;
localparam INT15 = 8'd143;
localparam INT16 = 8'd144;
localparam INT17 = 8'd145;
localparam INT18 = 8'd146;
localparam INT19 = 8'd147;
localparam INT20 = 8'd148;
localparam INT21 = 8'd149;
localparam INT22 = 8'd150;
localparam INT23 = 8'd151;
localparam INT24 = 8'd152;
localparam INT25 = 8'd153;
localparam INT26 = 8'd154;
localparam INT27 = 8'd155;
localparam INT28 = 8'd156;
localparam INT29 = 8'd157;
localparam INT30 = 8'd158;
localparam INT31 = 8'd159;
localparam INT32 = 8'd160;
localparam INT33 = 8'd161;
localparam INT34 = 8'd162;
localparam INT35 = 8'd163;
localparam INT36 = 8'd164;
localparam INT37 = 8'd165;
localparam INT38 = 8'd166;
localparam INT39 = 8'd167;
localparam INT40 = 8'd168;
localparam INT41 = 8'd169;
localparam INT42 = 8'd170;
localparam INT43 = 8'd171;
localparam INT44 = 8'd172;
localparam INT45 = 8'd173;
localparam INT46 = 8'd174;
localparam INT47 = 8'd175;
localparam INT48 = 8'd176;
localparam INT49 = 8'd177;
localparam INT50 = 8'd178;
localparam INT51 = 8'd179;
localparam INT52 = 8'd180;
localparam INT53 = 8'd181;
localparam INT54 = 8'd182;
localparam INT55 = 8'd183;
localparam INT56 = 8'd184;
localparam INT57 = 8'd185;
localparam INT58 = 8'd186;
localparam INT59 = 8'd187;
localparam INT60 = 8'd188;
localparam INT61 = 8'd189;
localparam INT62 = 8'd190;
localparam INT63 = 8'd191;
localparam INT64 = 8'd192;

// NEG_INT1 to NEG_INT16
localparam NEG_INT1 = 8'd193;
localparam NEG_INT2 = 8'd194;
localparam NEG_INT3 = 8'd195;
localparam NEG_INT4 = 8'd196;
localparam NEG_INT5 = 8'd197;
localparam NEG_INT6 = 8'd198;
localparam NEG_INT7 = 8'd199;
localparam NEG_INT8 = 8'd200;
localparam NEG_INT9 = 8'd201;
localparam NEG_INT10 = 8'd202;
localparam NEG_INT11 = 8'd203;
localparam NEG_INT12 = 8'd204;
localparam NEG_INT13 = 8'd205;
localparam NEG_INT14 = 8'd206;
localparam NEG_INT15 = 8'd207;
localparam NEG_INT16 = 8'd208;

localparam DPP8 = 8'd233;
localparam DPP8FI = 8'd233;
localparam SHARED_BASE = 8'd235;
localparam SHARED_LIMIT = 8'd236;
localparam PRIVATE_BASE = 8'd237;
localparam PRIVATE_LIMIT = 8'd238;
localparam POPS_EXITING_WAVE_ID = 8'd239;
localparam FLOAT_0_5 = 8'd240;
localparam FLOAT_NEG_0_5 = 8'd241;
localparam FLOAT_1_0 = 8'd242;
localparam FLOAT_NEG_1_0 = 8'd243;
localparam FLOAT_2_0 = 8'd244;
localparam FLOAT_NEG_2_0 = 8'd245;
localparam FLOAT_4_0 = 8'd246;
localparam FLOAT_NEG_4_0 = 8'd247;
localparam INV_TWO_PI = 8'd248;
localparam SDWA = 8'd249;
localparam RESERVED_249 = 8'd249;  // Reserved values 249-250
localparam DPP16 = 8'd250;
localparam RESERVED_250 = 8'd250;
localparam VCCZ = 8'd251;
localparam EXECZ = 8'd252;
localparam SCC = 8'd253;
localparam RESERVED_254 = 8'd254;
localparam LITERAL_CONSTANT = 8'd255;

// Vector Source Localparams
localparam S_VGPR0    = 9'd256;
localparam S_VGPR1    = 9'd257;
localparam S_VGPR2    = 9'd258;
localparam S_VGPR3    = 9'd259;
localparam S_VGPR4    = 9'd260;
localparam S_VGPR5    = 9'd261;
localparam S_VGPR6    = 9'd262;
localparam S_VGPR7    = 9'd263;
localparam S_VGPR8    = 9'd264;
localparam S_VGPR9    = 9'd265;
localparam S_VGPR10   = 9'd266;
localparam S_VGPR11   = 9'd267;
localparam S_VGPR12   = 9'd268;
localparam S_VGPR13   = 9'd269;
localparam S_VGPR14   = 9'd270;
localparam S_VGPR15   = 9'd271;
localparam S_VGPR16   = 9'd272;
localparam S_VGPR17   = 9'd273;
localparam S_VGPR18   = 9'd274;
localparam S_VGPR19   = 9'd275;
localparam S_VGPR20   = 9'd276;
localparam S_VGPR21   = 9'd277;
localparam S_VGPR22   = 9'd278;
localparam S_VGPR23   = 9'd279;
localparam S_VGPR24   = 9'd280;
localparam S_VGPR25   = 9'd281;
localparam S_VGPR26   = 9'd282;
localparam S_VGPR27   = 9'd283;
localparam S_VGPR28   = 9'd284;
localparam S_VGPR29   = 9'd285;
localparam S_VGPR30   = 9'd286;
localparam S_VGPR31   = 9'd287;
localparam S_VGPR32   = 9'd288;
localparam S_VGPR33   = 9'd289;
localparam S_VGPR34   = 9'd290;
localparam S_VGPR35   = 9'd291;
localparam S_VGPR36   = 9'd292;
localparam S_VGPR37   = 9'd293;
localparam S_VGPR38   = 9'd294;
localparam S_VGPR39   = 9'd295;
localparam S_VGPR40   = 9'd296;
localparam S_VGPR41   = 9'd297;
localparam S_VGPR42   = 9'd298;
localparam S_VGPR43   = 9'd299;
localparam S_VGPR44   = 9'd300;
localparam S_VGPR45   = 9'd301;
localparam S_VGPR46   = 9'd302;
localparam S_VGPR47   = 9'd303;
localparam S_VGPR48   = 9'd304;
localparam S_VGPR49   = 9'd305;
localparam S_VGPR50   = 9'd306;
localparam S_VGPR51   = 9'd307;
localparam S_VGPR52   = 9'd308;
localparam S_VGPR53   = 9'd309;
localparam S_VGPR54   = 9'd310;
localparam S_VGPR55   = 9'd311;
localparam S_VGPR56   = 9'd312;
localparam S_VGPR57   = 9'd313;
localparam S_VGPR58   = 9'd314;
localparam S_VGPR59   = 9'd315;
localparam S_VGPR60   = 9'd316;
localparam S_VGPR61   = 9'd317;
localparam S_VGPR62   = 9'd318;
localparam S_VGPR63   = 9'd319;
localparam S_VGPR64   = 9'd320;
localparam S_VGPR65   = 9'd321;
localparam S_VGPR66   = 9'd322;
localparam S_VGPR67   = 9'd323;
localparam S_VGPR68   = 9'd324;
localparam S_VGPR69   = 9'd325;
localparam S_VGPR70   = 9'd326;
localparam S_VGPR71   = 9'd327;
localparam S_VGPR72   = 9'd328;
localparam S_VGPR73   = 9'd329;
localparam S_VGPR74   = 9'd330;
localparam S_VGPR75   = 9'd331;
localparam S_VGPR76   = 9'd332;
localparam S_VGPR77   = 9'd333;
localparam S_VGPR78   = 9'd334;
localparam S_VGPR79   = 9'd335;
localparam S_VGPR80   = 9'd336;
localparam S_VGPR81   = 9'd337;
localparam S_VGPR82   = 9'd338;
localparam S_VGPR83   = 9'd339;
localparam S_VGPR84   = 9'd340;
localparam S_VGPR85   = 9'd341;
localparam S_VGPR86   = 9'd342;
localparam S_VGPR87   = 9'd343;
localparam S_VGPR88   = 9'd344;
localparam S_VGPR89   = 9'd345;
localparam S_VGPR90   = 9'd346;
localparam S_VGPR91   = 9'd347;
localparam S_VGPR92   = 9'd348;
localparam S_VGPR93   = 9'd349;
localparam S_VGPR94   = 9'd350;
localparam S_VGPR95   = 9'd351;
localparam S_VGPR96   = 9'd352;
localparam S_VGPR97   = 9'd353;
localparam S_VGPR98   = 9'd354;
localparam S_VGPR99   = 9'd355;
localparam S_VGPR100  = 9'd356;
localparam S_VGPR101  = 9'd357;
localparam S_VGPR102  = 9'd358;
localparam S_VGPR103  = 9'd359;
localparam S_VGPR104  = 9'd360;
localparam S_VGPR105  = 9'd361;
localparam S_VGPR106  = 9'd362;
localparam S_VGPR107  = 9'd363;
localparam S_VGPR108  = 9'd364;
localparam S_VGPR109  = 9'd365;
localparam S_VGPR110  = 9'd366;
localparam S_VGPR111  = 9'd367;
localparam S_VGPR112  = 9'd368;
localparam S_VGPR113  = 9'd369;
localparam S_VGPR114  = 9'd370;
localparam S_VGPR115  = 9'd371;
localparam S_VGPR116  = 9'd372;
localparam S_VGPR117  = 9'd373;
localparam S_VGPR118  = 9'd374;
localparam S_VGPR119  = 9'd375;
localparam S_VGPR120  = 9'd376;
localparam S_VGPR121  = 9'd377;
localparam S_VGPR122  = 9'd378;
localparam S_VGPR123  = 9'd379;
localparam S_VGPR124  = 9'd380;
localparam S_VGPR125  = 9'd381;
localparam S_VGPR126  = 9'd382;
localparam S_VGPR127  = 9'd383;
localparam S_VGPR128  = 9'd384;
localparam S_VGPR129  = 9'd385;
localparam S_VGPR130  = 9'd386;
localparam S_VGPR131  = 9'd387;
localparam S_VGPR132  = 9'd388;
localparam S_VGPR133  = 9'd389;
localparam S_VGPR134  = 9'd390;
localparam S_VGPR135  = 9'd391;
localparam S_VGPR136  = 9'd392;
localparam S_VGPR137  = 9'd393;
localparam S_VGPR138  = 9'd394;
localparam S_VGPR139  = 9'd395;
localparam S_VGPR140  = 9'd396;
localparam S_VGPR141  = 9'd397;
localparam S_VGPR142  = 9'd398;
localparam S_VGPR143  = 9'd399;
localparam S_VGPR144  = 9'd400;
localparam S_VGPR145  = 9'd401;
localparam S_VGPR146  = 9'd402;
localparam S_VGPR147  = 9'd403;
localparam S_VGPR148  = 9'd404;
localparam S_VGPR149  = 9'd405;
localparam S_VGPR150  = 9'd406;
localparam S_VGPR151  = 9'd407;
localparam S_VGPR152  = 9'd408;
localparam S_VGPR153  = 9'd409;
localparam S_VGPR154  = 9'd410;
localparam S_VGPR155  = 9'd411;
localparam S_VGPR156  = 9'd412;
localparam S_VGPR157  = 9'd413;
localparam S_VGPR158  = 9'd414;
localparam S_VGPR159  = 9'd415;
localparam S_VGPR160  = 9'd416;
localparam S_VGPR161  = 9'd417;
localparam S_VGPR162  = 9'd418;
localparam S_VGPR163  = 9'd419;
localparam S_VGPR164  = 9'd420;
localparam S_VGPR165  = 9'd421;
localparam S_VGPR166  = 9'd422;
localparam S_VGPR167  = 9'd423;
localparam S_VGPR168  = 9'd424;
localparam S_VGPR169  = 9'd425;
localparam S_VGPR170  = 9'd426;
localparam S_VGPR171  = 9'd427;
localparam S_VGPR172  = 9'd428;
localparam S_VGPR173  = 9'd429;
localparam S_VGPR174  = 9'd430;
localparam S_VGPR175  = 9'd431;
localparam S_VGPR176  = 9'd432;
localparam S_VGPR177  = 9'd433;
localparam S_VGPR178  = 9'd434;
localparam S_VGPR179  = 9'd435;
localparam S_VGPR180  = 9'd436;
localparam S_VGPR181  = 9'd437;
localparam S_VGPR182  = 9'd438;
localparam S_VGPR183  = 9'd439;
localparam S_VGPR184  = 9'd440;
localparam S_VGPR185  = 9'd441;
localparam S_VGPR186  = 9'd442;
localparam S_VGPR187  = 9'd443;
localparam S_VGPR188  = 9'd444;
localparam S_VGPR189  = 9'd445;
localparam S_VGPR190  = 9'd446;
localparam S_VGPR191  = 9'd447;
localparam S_VGPR192  = 9'd448;
localparam S_VGPR193  = 9'd449;
localparam S_VGPR194  = 9'd450;
localparam S_VGPR195  = 9'd451;
localparam S_VGPR196  = 9'd452;
localparam S_VGPR197  = 9'd453;
localparam S_VGPR198  = 9'd454;
localparam S_VGPR199  = 9'd455;
localparam S_VGPR200  = 9'd456;
localparam S_VGPR201  = 9'd457;
localparam S_VGPR202  = 9'd458;
localparam S_VGPR203  = 9'd459;
localparam S_VGPR204  = 9'd460;
localparam S_VGPR205  = 9'd461;
localparam S_VGPR206  = 9'd462;
localparam S_VGPR207  = 9'd463;
localparam S_VGPR208  = 9'd464;
localparam S_VGPR209  = 9'd465;
localparam S_VGPR210  = 9'd466;
localparam S_VGPR211  = 9'd467;
localparam S_VGPR212  = 9'd468;
localparam S_VGPR213  = 9'd469;
localparam S_VGPR214  = 9'd470;
localparam S_VGPR215  = 9'd471;
localparam S_VGPR216  = 9'd472;
localparam S_VGPR217  = 9'd473;
localparam S_VGPR218  = 9'd474;
localparam S_VGPR219  = 9'd475;
localparam S_VGPR220  = 9'd476;
localparam S_VGPR221  = 9'd477;
localparam S_VGPR222  = 9'd478;
localparam S_VGPR223  = 9'd479;
localparam S_VGPR224  = 9'd480;
localparam S_VGPR225  = 9'd481;
localparam S_VGPR226  = 9'd482;
localparam S_VGPR227  = 9'd483;
localparam S_VGPR228  = 9'd484;
localparam S_VGPR229  = 9'd485;
localparam S_VGPR230  = 9'd486;
localparam S_VGPR231  = 9'd487;
localparam S_VGPR232  = 9'd488;
localparam S_VGPR233  = 9'd489;
localparam S_VGPR234  = 9'd490;
localparam S_VGPR235  = 9'd491;
localparam S_VGPR236  = 9'd492;
localparam S_VGPR237  = 9'd493;
localparam S_VGPR238  = 9'd494;
localparam S_VGPR239  = 9'd495;
localparam S_VGPR240  = 9'd496;
localparam S_VGPR241  = 9'd497;
localparam S_VGPR242  = 9'd498;
localparam S_VGPR243  = 9'd499;
localparam S_VGPR244  = 9'd500;
localparam S_VGPR245  = 9'd501;
localparam S_VGPR246  = 9'd502;
localparam S_VGPR247  = 9'd503;
localparam S_VGPR248  = 9'd504;
localparam S_VGPR249  = 9'd505;
localparam S_VGPR250  = 9'd506;
localparam S_VGPR251  = 9'd507;
localparam S_VGPR252  = 9'd508;
localparam S_VGPR253  = 9'd509;
localparam S_VGPR254  = 9'd510;
localparam S_VGPR255  = 9'd511;

// Vector VSource Localparams
localparam VGPR0    = 8'd0;
localparam VGPR1    = 8'd1;
localparam VGPR2    = 8'd2;
localparam VGPR3    = 8'd3;
localparam VGPR4    = 8'd4;
localparam VGPR5    = 8'd5;
localparam VGPR6    = 8'd6;
localparam VGPR7    = 8'd7;
localparam VGPR8    = 8'd8;
localparam VGPR9    = 8'd9;
localparam VGPR10   = 8'd10;
localparam VGPR11   = 8'd11;
localparam VGPR12   = 8'd12;
localparam VGPR13   = 8'd13;
localparam VGPR14   = 8'd14;
localparam VGPR15   = 8'd15;
localparam VGPR16   = 8'd16;
localparam VGPR17   = 8'd17;
localparam VGPR18   = 8'd18;
localparam VGPR19   = 8'd19;
localparam VGPR20   = 8'd20;
localparam VGPR21   = 8'd21;
localparam VGPR22   = 8'd22;
localparam VGPR23   = 8'd23;
localparam VGPR24   = 8'd24;
localparam VGPR25   = 8'd25;
localparam VGPR26   = 8'd26;
localparam VGPR27   = 8'd27;
localparam VGPR28   = 8'd28;
localparam VGPR29   = 8'd29;
localparam VGPR30   = 8'd30;
localparam VGPR31   = 8'd31;
localparam VGPR32   = 8'd32;
localparam VGPR33   = 8'd33;
localparam VGPR34   = 8'd34;
localparam VGPR35   = 8'd35;
localparam VGPR36   = 8'd36;
localparam VGPR37   = 8'd37;
localparam VGPR38   = 8'd38;
localparam VGPR39   = 8'd39;
localparam VGPR40   = 8'd40;
localparam VGPR41   = 8'd41;
localparam VGPR42   = 8'd42;
localparam VGPR43   = 8'd43;
localparam VGPR44   = 8'd44;
localparam VGPR45   = 8'd45;
localparam VGPR46   = 8'd46;
localparam VGPR47   = 8'd47;
localparam VGPR48   = 8'd48;
localparam VGPR49   = 8'd49;
localparam VGPR50   = 8'd50;
localparam VGPR51   = 8'd51;
localparam VGPR52   = 8'd52;
localparam VGPR53   = 8'd53;
localparam VGPR54   = 8'd54;
localparam VGPR55   = 8'd55;
localparam VGPR56   = 8'd56;
localparam VGPR57   = 8'd57;
localparam VGPR58   = 8'd58;
localparam VGPR59   = 8'd59;
localparam VGPR60   = 8'd60;
localparam VGPR61   = 8'd61;
localparam VGPR62   = 8'd62;
localparam VGPR63   = 8'd63;
localparam VGPR64   = 8'd64;
localparam VGPR65   = 8'd65;
localparam VGPR66   = 8'd66;
localparam VGPR67   = 8'd67;
localparam VGPR68   = 8'd68;
localparam VGPR69   = 8'd69;
localparam VGPR70   = 8'd70;
localparam VGPR71   = 8'd71;
localparam VGPR72   = 8'd72;
localparam VGPR73   = 8'd73;
localparam VGPR74   = 8'd74;
localparam VGPR75   = 8'd75;
localparam VGPR76   = 8'd76;
localparam VGPR77   = 8'd77;
localparam VGPR78   = 8'd78;
localparam VGPR79   = 8'd79;
localparam VGPR80   = 8'd80;
localparam VGPR81   = 8'd81;
localparam VGPR82   = 8'd82;
localparam VGPR83   = 8'd83;
localparam VGPR84   = 8'd84;
localparam VGPR85   = 8'd85;
localparam VGPR86   = 8'd86;
localparam VGPR87   = 8'd87;
localparam VGPR88   = 8'd88;
localparam VGPR89   = 8'd89;
localparam VGPR90   = 8'd90;
localparam VGPR91   = 8'd91;
localparam VGPR92   = 8'd92;
localparam VGPR93   = 8'd93;
localparam VGPR94   = 8'd94;
localparam VGPR95   = 8'd95;
localparam VGPR96   = 8'd96;
localparam VGPR97   = 8'd97;
localparam VGPR98   = 8'd98;
localparam VGPR99   = 8'd99;
localparam VGPR100  = 8'd100;
localparam VGPR101  = 8'd101;
localparam VGPR102  = 8'd102;
localparam VGPR103  = 8'd103;
localparam VGPR104  = 8'd104;
localparam VGPR105  = 8'd105;
localparam VGPR106  = 8'd106;
localparam VGPR107  = 8'd107;
localparam VGPR108  = 8'd108;
localparam VGPR109  = 8'd109;
localparam VGPR110  = 8'd110;
localparam VGPR111  = 8'd111;
localparam VGPR112  = 8'd112;
localparam VGPR113  = 8'd113;
localparam VGPR114  = 8'd114;
localparam VGPR115  = 8'd115;
localparam VGPR116  = 8'd116;
localparam VGPR117  = 8'd117;
localparam VGPR118  = 8'd118;
localparam VGPR119  = 8'd119;
localparam VGPR120  = 8'd120;
localparam VGPR121  = 8'd121;
localparam VGPR122  = 8'd122;
localparam VGPR123  = 8'd123;
localparam VGPR124  = 8'd124;
localparam VGPR125  = 8'd125;
localparam VGPR126  = 8'd126;
localparam VGPR127  = 8'd127;
localparam VGPR128  = 8'd128;
localparam VGPR129  = 8'd129;
localparam VGPR130  = 8'd130;
localparam VGPR131  = 8'd131;
localparam VGPR132  = 8'd132;
localparam VGPR133  = 8'd133;
localparam VGPR134  = 8'd134;
localparam VGPR135  = 8'd135;
localparam VGPR136  = 8'd136;
localparam VGPR137  = 8'd137;
localparam VGPR138  = 8'd138;
localparam VGPR139  = 8'd139;
localparam VGPR140  = 8'd140;
localparam VGPR141  = 8'd141;
localparam VGPR142  = 8'd142;
localparam VGPR143  = 8'd143;
localparam VGPR144  = 8'd144;
localparam VGPR145  = 8'd145;
localparam VGPR146  = 8'd146;
localparam VGPR147  = 8'd147;
localparam VGPR148  = 8'd148;
localparam VGPR149  = 8'd149;
localparam VGPR150  = 8'd150;
localparam VGPR151  = 8'd151;
localparam VGPR152  = 8'd152;
localparam VGPR153  = 8'd153;
localparam VGPR154  = 8'd154;
localparam VGPR155  = 8'd155;
localparam VGPR156  = 8'd156;
localparam VGPR157  = 8'd157;
localparam VGPR158  = 8'd158;
localparam VGPR159  = 8'd159;
localparam VGPR160  = 8'd160;
localparam VGPR161  = 8'd161;
localparam VGPR162  = 8'd162;
localparam VGPR163  = 8'd163;
localparam VGPR164  = 8'd164;
localparam VGPR165  = 8'd165;
localparam VGPR166  = 8'd166;
localparam VGPR167  = 8'd167;
localparam VGPR168  = 8'd168;
localparam VGPR169  = 8'd169;
localparam VGPR170  = 8'd170;
localparam VGPR171  = 8'd171;
localparam VGPR172  = 8'd172;
localparam VGPR173  = 8'd173;
localparam VGPR174  = 8'd174;
localparam VGPR175  = 8'd175;
localparam VGPR176  = 8'd176;
localparam VGPR177  = 8'd177;
localparam VGPR178  = 8'd178;
localparam VGPR179  = 8'd179;
localparam VGPR180  = 8'd180;
localparam VGPR181  = 8'd181;
localparam VGPR182  = 8'd182;
localparam VGPR183  = 8'd183;
localparam VGPR184  = 8'd184;
localparam VGPR185  = 8'd185;
localparam VGPR186  = 8'd186;
localparam VGPR187  = 8'd187;
localparam VGPR188  = 8'd188;
localparam VGPR189  = 8'd189;
localparam VGPR190  = 8'd190;
localparam VGPR191  = 8'd191;
localparam VGPR192  = 8'd192;
localparam VGPR193  = 8'd193;
localparam VGPR194  = 8'd194;
localparam VGPR195  = 8'd195;
localparam VGPR196  = 8'd196;
localparam VGPR197  = 8'd197;
localparam VGPR198  = 8'd198;
localparam VGPR199  = 8'd199;
localparam VGPR200  = 8'd200;
localparam VGPR201  = 8'd201;
localparam VGPR202  = 8'd202;
localparam VGPR203  = 8'd203;
localparam VGPR204  = 8'd204;
localparam VGPR205  = 8'd205;
localparam VGPR206  = 8'd206;
localparam VGPR207  = 8'd207;
localparam VGPR208  = 8'd208;
localparam VGPR209  = 8'd209;
localparam VGPR210  = 8'd210;
localparam VGPR211  = 8'd211;
localparam VGPR212  = 8'd212;
localparam VGPR213  = 8'd213;
localparam VGPR214  = 8'd214;
localparam VGPR215  = 8'd215;
localparam VGPR216  = 8'd216;
localparam VGPR217  = 8'd217;
localparam VGPR218  = 8'd218;
localparam VGPR219  = 8'd219;
localparam VGPR220  = 8'd220;
localparam VGPR221  = 8'd221;
localparam VGPR222  = 8'd222;
localparam VGPR223  = 8'd223;
localparam VGPR224  = 8'd224;
localparam VGPR225  = 8'd225;
localparam VGPR226  = 8'd226;
localparam VGPR227  = 8'd227;
localparam VGPR228  = 8'd228;
localparam VGPR229  = 8'd229;
localparam VGPR230  = 8'd230;
localparam VGPR231  = 8'd231;
localparam VGPR232  = 8'd232;
localparam VGPR233  = 8'd233;
localparam VGPR234  = 8'd234;
localparam VGPR235  = 8'd235;
localparam VGPR236  = 8'd236;
localparam VGPR237  = 8'd237;
localparam VGPR238  = 8'd238;
localparam VGPR239  = 8'd239;
localparam VGPR240  = 8'd240;
localparam VGPR241  = 8'd241;
localparam VGPR242  = 8'd242;
localparam VGPR243  = 8'd243;
localparam VGPR244  = 8'd244;
localparam VGPR245  = 8'd245;
localparam VGPR246  = 8'd246;
localparam VGPR247  = 8'd247;
localparam VGPR248  = 8'd248;
localparam VGPR249  = 8'd249;
localparam VGPR250  = 8'd250;
localparam VGPR251  = 8'd251;
localparam VGPR252  = 8'd252;
localparam VGPR253  = 8'd253;
localparam VGPR254  = 8'd254;
localparam VGPR255  = 8'd255;

endpackage
