package arithmetic_pkg;

typedef enum {
    LSHFTL,
    LSHFTR,
    ASHFTR,
    AND,
    XOR,
    OR,
    S_LT,
    S_GT,
    U_LT,
    U_GT,
    EQ,
    MAX3
} logic_op_t;

endpackage
