`timescale 1ps/1ps

package flat_op_pkg; 

    localparam GLOBAL_LOAD_DWORD    = 7'd12;
    localparam GLOBAL_LOAD_DWORDX2  = 7'd13;

    localparam GLOBAL_STORE_DWORD   = 7'd28;

endpackage
