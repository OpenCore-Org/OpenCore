`timescale 1ps/1ps

package scalar_op_pkg; 

    // SOP2 instruction opcodes
    localparam SOP2_ADD_U32             = 8'd0;
    localparam SOP2_SUB_U32             = 8'd1;
    localparam SOP2_ADD_I32             = 8'd2;
    localparam SOP2_SUB_I32             = 8'd3;
    localparam SOP2_ADDC_U32            = 8'd4;
    localparam SOP2_SUBB_U32            = 8'd5;
    localparam SOP2_MIN_I32             = 8'd6;
    localparam SOP2_MIN_U32             = 8'd7;
    localparam SOP2_MAX_I32             = 8'd8;
    localparam SOP2_MAX_U32             = 8'd9;
    localparam SOP2_CSELECT_B32         = 8'd10;
    localparam SOP2_CSELECT_B64         = 8'd11;
    localparam SOP2_AND_B32             = 8'd14;
    localparam SOP2_AND_B64             = 8'd15;
    localparam SOP2_OR_B32              = 8'd16;
    localparam SOP2_OR_B64              = 8'd17;
    localparam SOP2_XOR_B32             = 8'd18;
    localparam SOP2_XOR_B64             = 8'd19;
    localparam SOP2_ANDN2_B32           = 8'd20;
    localparam SOP2_ANDN2_B64           = 8'd21;
    localparam SOP2_ORN2_B32            = 8'd22;
    localparam SOP2_ORN2_B64            = 8'd23;
    localparam SOP2_NAND_B32            = 8'd24;
    localparam SOP2_NAND_B64            = 8'd25;
    localparam SOP2_NOR_B32             = 8'd26;
    localparam SOP2_NOR_B64             = 8'd27;
    localparam SOP2_XNOR_B32            = 8'd28;
    localparam SOP2_XNOR_B64            = 8'd29;
    localparam SOP2_LSHL_B32            = 8'd30;
    localparam SOP2_LSHL_B64            = 8'd31;
    localparam SOP2_LSHR_B32            = 8'd32;
    localparam SOP2_LSHR_B64            = 8'd33;
    localparam SOP2_ASHR_I32            = 8'd34;
    localparam SOP2_ASHR_I64            = 8'd35;
    localparam SOP2_BFM_B32             = 8'd36;
    localparam SOP2_BFM_B64             = 8'd37;
    localparam SOP2_MUL_I32             = 8'd38;
    localparam SOP2_BFE_U32             = 8'd39;
    localparam SOP2_BFE_I32             = 8'd40;
    localparam SOP2_BFE_U64             = 8'd41;
    localparam SOP2_BFE_I64             = 8'd42;
    localparam SOP2_ABSDIFF_I32         = 8'd44;
    localparam SOP2_LSHL1_ADD_U32       = 8'd46;
    localparam SOP2_LSHL2_ADD_U32       = 8'd47;
    localparam SOP2_LSHL3_ADD_U32       = 8'd48;
    localparam SOP2_LSHL4_ADD_U32       = 8'd49;
    localparam SOP2_PACK_LL_B32_B16     = 8'd50;
    localparam SOP2_PACK_LH_B32_B16     = 8'd51;
    localparam SOP2_PACK_HH_B32_B16     = 8'd52;
    localparam SOP2_MUL_HI_U32          = 8'd53;
    localparam SOP2_MUL_HI_I32          = 8'd54;

    // SOP1 instruction opcodes
    localparam SOP1_MOV_B32                = 8'd3;
    localparam SOP1_MOV_B64                = 8'd4;
    localparam SOP1_CMOV_B32               = 8'd5;
    localparam SOP1_CMOV_B64               = 8'd6;
    localparam SOP1_NOT_B32                = 8'd7;
    localparam SOP1_NOT_B64                = 8'd8;
    localparam SOP1_WQM_B32                = 8'd9;
    localparam SOP1_WQM_B64                = 8'd10;
    localparam SOP1_BREV_B32               = 8'd11;
    localparam SOP1_BREV_B64               = 8'd12;
    localparam SOP1_BCNT0_I32_B32          = 8'd13;
    localparam SOP1_BCNT0_I32_B64          = 8'd14;
    localparam SOP1_BCNT1_I32_B32          = 8'd15;
    localparam SOP1_BCNT1_I32_B64          = 8'd16;
    localparam SOP1_FF0_I32_B32            = 8'd17;
    localparam SOP1_FF0_I32_B64            = 8'd18;
    localparam SOP1_FF1_I32_B32            = 8'd19;
    localparam SOP1_FF1_I32_B64            = 8'd20;
    localparam SOP1_FLBIT_I32_B32          = 8'd21;
    localparam SOP1_FLBIT_I32_B64          = 8'd22;
    localparam SOP1_FLBIT_I32              = 8'd23;
    localparam SOP1_FLBIT_I32_I64          = 8'd24;
    localparam SOP1_SEXT_I32_I8            = 8'd25;
    localparam SOP1_SEXT_I32_I16           = 8'd26;
    localparam SOP1_BITSET0_B32            = 8'd27;
    localparam SOP1_BITSET0_B64            = 8'd28;
    localparam SOP1_BITSET1_B32            = 8'd29;
    localparam SOP1_BITSET1_B64            = 8'd30;
    localparam SOP1_GETPC_B64              = 8'd31;
    localparam SOP1_SETPC_B64              = 8'd32;
    localparam SOP1_SWAPPC_B64             = 8'd33;
    localparam SOP1_RFE_B64                = 8'd34;
    localparam SOP1_AND_SAVEEXEC_B64       = 8'd36;
    localparam SOP1_OR_SAVEEXEC_B64        = 8'd37;
    localparam SOP1_XOR_SAVEEXEC_B64       = 8'd38;
    localparam SOP1_ANDN2_SAVEEXEC_B64     = 8'd39;
    localparam SOP1_ORN2_SAVEEXEC_B64      = 8'd40;
    localparam SOP1_NAND_SAVEEXEC_B64      = 8'd41;
    localparam SOP1_NOR_SAVEEXEC_B64       = 8'd42;
    localparam SOP1_XNOR_SAVEEXEC_B64      = 8'd43;
    localparam SOP1_QUADMASK_B32           = 8'd44;
    localparam SOP1_QUADMASK_B64           = 8'd45;
    localparam SOP1_MOVRELS_B32            = 8'd46;
    localparam SOP1_MOVRELS_B64            = 8'd47;
    localparam SOP1_MOVRELD_B32            = 8'd48;
    localparam SOP1_MOVRELD_B64            = 8'd49;
    localparam SOP1_ABS_I32                = 8'd52;
    localparam SOP1_ANDN1_SAVEEXEC_B64     = 8'd55;
    localparam SOP1_ORN1_SAVEEXEC_B64      = 8'd56;
    localparam SOP1_ANDN1_WREXEC_B64       = 8'd57;
    localparam SOP1_ANDN2_WREXEC_B64       = 8'd58;
    localparam SOP1_BITREPLICATE_B64_B32   = 8'd59;
    localparam SOP1_AND_SAVEEXEC_B32       = 8'd60;
    localparam SOP1_OR_SAVEEXEC_B32        = 8'd61;
    localparam SOP1_XOR_SAVEEXEC_B32       = 8'd62;
    localparam SOP1_ANDN2_SAVEEXEC_B32     = 8'd63;
    localparam SOP1_ORN2_SAVEEXEC_B32      = 8'd64;
    localparam SOP1_NAND_SAVEEXEC_B32      = 8'd65;
    localparam SOP1_NOR_SAVEEXEC_B32       = 8'd66;
    localparam SOP1_XNOR_SAVEEXEC_B32      = 8'd67;
    localparam SOP1_ANDN1_SAVEEXEC_B32     = 8'd68;
    localparam SOP1_ORN1_SAVEEXEC_B32      = 8'd69;
    localparam SOP1_ANDN1_WREXEC_B32       = 8'd70;
    localparam SOP1_ANDN2_WREXEC_B32       = 8'd71;
    localparam SOP1_MOVRELSD_2_B32         = 8'd73;

    // SOPK instruction opcodes
    localparam SOPK_MOVK_I32               = 8'd0;
    localparam SOPK_VERSION                = 8'd1;
    localparam SOPK_CMOVK_I32              = 8'd2;
    localparam SOPK_CMPK_EQ_I32            = 8'd3;
    localparam SOPK_CMPK_LG_I32            = 8'd4;
    localparam SOPK_CMPK_GT_I32            = 8'd5;
    localparam SOPK_CMPK_GE_I32            = 8'd6;
    localparam SOPK_CMPK_LT_I32            = 8'd7;
    localparam SOPK_CMPK_LE_I32            = 8'd8;
    localparam SOPK_CMPK_EQ_U32            = 8'd9;
    localparam SOPK_CMPK_LG_U32            = 8'd10;
    localparam SOPK_CMPK_GT_U32            = 8'd11;
    localparam SOPK_CMPK_GE_U32            = 8'd12;
    localparam SOPK_CMPK_LT_U32            = 8'd13;
    localparam SOPK_CMPK_LE_U32            = 8'd14;
    localparam SOPK_ADDK_I32               = 8'd15;
    localparam SOPK_MULK_I32               = 8'd16;
    localparam SOPK_GETREG_B32             = 8'd18;
    localparam SOPK_SETREG_B32             = 8'd19;
    localparam SOPK_SETREG_IMM32_B32       = 8'd21;
    localparam SOPK_CALL_B64               = 8'd22;
    localparam SOPK_WAITCNT_VSCNT          = 8'd23;
    localparam SOPK_WAITCNT_VMCNT          = 8'd24;
    localparam SOPK_WAITCNT_EXPCNT         = 8'd25;
    localparam SOPK_WAITCNT_LGKMCNT        = 8'd26;
    localparam SOPK_SUBVECTOR_LOOP_BEGIN   = 8'd27;
    localparam SOPK_SUBVECTOR_LOOP_END     = 8'd28;

    // SOPC instruction opcodes
    localparam SOPC_CMP_EQ_I32             = 8'd0;
    localparam SOPC_CMP_LG_I32             = 8'd1;
    localparam SOPC_CMP_GT_I32             = 8'd2;
    localparam SOPC_CMP_GE_I32             = 8'd3;
    localparam SOPC_CMP_LT_I32             = 8'd4;
    localparam SOPC_CMP_LE_I32             = 8'd5;
    localparam SOPC_CMP_EQ_U32             = 8'd6;
    localparam SOPC_CMP_LG_U32             = 8'd7;
    localparam SOPC_CMP_GT_U32             = 8'd8;
    localparam SOPC_CMP_GE_U32             = 8'd9;
    localparam SOPC_CMP_LT_U32             = 8'd10;
    localparam SOPC_CMP_LE_U32             = 8'd11;
    localparam SOPC_BITCMP0_B32            = 8'd12;
    localparam SOPC_BITCMP1_B32            = 8'd13;
    localparam SOPC_BITCMP0_B64            = 8'd14;
    localparam SOPC_BITCMP1_B64            = 8'd15;
    localparam SOPC_CMP_EQ_U64             = 8'd18;
    localparam SOPC_CMP_LG_U64             = 8'd19;

    // SOPP instruction opcodes
    localparam SOPP_NOP                        = 8'd0;
    localparam SOPP_ENDPGM                     = 8'd1;
    localparam SOPP_BRANCH                     = 8'd2;
    localparam SOPP_WAKEUP                     = 8'd3;
    localparam SOPP_CBRANCH_SCC0               = 8'd4;
    localparam SOPP_CBRANCH_SCC1               = 8'd5;
    localparam SOPP_CBRANCH_VCCZ               = 8'd6;
    localparam SOPP_CBRANCH_VCCNZ              = 8'd7;
    localparam SOPP_CBRANCH_EXECZ              = 8'd8;
    localparam SOPP_CBRANCH_EXECNZ             = 8'd9;
    localparam SOPP_BARRIER                    = 8'd10;
    localparam SOPP_SETKILL                    = 8'd11;
    localparam SOPP_WAITCNT                    = 8'd12;
    localparam SOPP_SETHALT                    = 8'd13;
    localparam SOPP_SLEEP                      = 8'd14;
    localparam SOPP_SETPRIO                    = 8'd15;
    localparam SOPP_SENDMSG                    = 8'd16;
    localparam SOPP_SENDMSGHALT                = 8'd17;
    localparam SOPP_TRAP                       = 8'd18;
    localparam SOPP_ICACHE_INV                 = 8'd19;
    localparam SOPP_INCPERFLEVEL               = 8'd20;
    localparam SOPP_DECPERFLEVEL               = 8'd21;
    localparam SOPP_TTRACEDATA                 = 8'd22;
    localparam SOPP_CBRANCH_CDBGSYS            = 8'd23;
    localparam SOPP_CBRANCH_CDBGUSER           = 8'd24;
    localparam SOPP_CBRANCH_CDBGSYS_OR_USER    = 8'd25;
    localparam SOPP_CBRANCH_CDBGSYS_AND_USER   = 8'd26;
    localparam SOPP_ENDPGM_SAVED               = 8'd27;
    localparam SOPP_ENDPGM_ORDERED_PS_DONE     = 8'd30;
    localparam SOPP_CODE_END                   = 8'd31;
    localparam SOPP_INST_PREFETCH              = 8'd32;
    localparam SOPP_CLAUSE                     = 8'd33;
    localparam SOPP_WAITCNT_DEPCTR             = 8'd35;
    localparam SOPP_ROUND_MODE                 = 8'd36;
    localparam SOPP_DENORM_MODE                = 8'd37;
    localparam SOPP_TTRACEDATA_IMM             = 8'd40;

endpackage
